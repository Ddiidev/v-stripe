module stripe

pub interface IStripe {
	secret_key string
}
