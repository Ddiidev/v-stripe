module stripe

pub struct Stripe {
pub:
	secret_key string
}
